endmodule
